endmodule
